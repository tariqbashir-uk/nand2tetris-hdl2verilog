module And(out, a, b);
    input a, b;
    output out;
    and(out, a, b);
endmodule