module Or(out, a, b);
    input a, b;
    output out;
    or(out, a, b);
endmodule