module Nand(out, a, b);
  input a, b;
  output out;
  nand (out, a, b);
endmodule