module Not(out, in);
    input in;
    output out;
    not (out, in);
endmodule